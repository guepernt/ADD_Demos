//ECE 6370
//David Zhang, 2213233

//This module counts to 100 based on the clk input. It is part of a nested loop that counts to a total
//of 50,000,000, at which point it will determine that 1 second has passed.

//For simulation purposes, this module will be set to a count of 3. The real number should be set
//back after simulation to be 7'b1100100, minus 1.
module countTo100(clk, rst, enable, counter_out);
	input clk, enable, rst;
	output counter_out;
	reg counter_out;

	reg [6:0] rollingCounter;
	wire counter_wire;
	parameter OFF = 0, ON = 1;
	reg State;
	countTo10 counter(clk, rst, enable, counter_wire);
	
	always @(posedge clk) begin
		if(rst == 1'b0) begin
			rollingCounter <= 7'b0000000;
			counter_out <= 1'b0;
			State <= OFF;
		end
		else
			case (State) 
				OFF: begin
					rollingCounter <= 0;
					counter_out <= 0;
					if (enable == 1'b1) begin
						State <= ON;
					end
				end

				ON: begin
					if (enable == 1'b1) begin
						if (counter_wire == 1'b1) begin
							if (rollingCounter == 7'b1100011) begin	//Set back after simulation
								counter_out <= 1'b1;
								rollingCounter <= 0;
							end
							else begin
								counter_out <= 1'b0;
								rollingCounter <= rollingCounter + 1'b1;
							end
						end
						else begin
							counter_out <= 1'b0;
						end
					end
					else begin
						State <= OFF;
					end
				end
		
				default: begin
					State <= OFF;
				end
			endcase
	end		
endmodule
